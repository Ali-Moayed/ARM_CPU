module test_bench(Din,clock,Aout,Bout,op);
output reg [63:0]Aout;
output reg [63:0]Bout;
output reg [3:0]op;
input clock;
input Din;
reg [131:0]c[7:0];
reg [63:0]d[7:0];

integer k = 0;
initial
begin
  c[0] = 132'b00111110000000000110000000000000000101010000000000011100100000111110110000000001100110011000000000000001101110000000100100010000000;
  c[1] = 132'b01010001111001111110000001111100000100000001100000011100100000000110110000010001100101000000000011110000100010011000100100000000001;
  c[2] = 132'b00001111100111000110000111000001110001100110110011000011110001000110000011110000010110011000011111001000010000000010100100010000010;
  c[3] = 132'b11100001110000000110001001001000000100010010010010000011100100110111011000100100001100110011000001100000001101110000000100100010110;
  c[4] = 132'b00100110011011000000000000100000010101000000010101001110010000101100000001100110011001100000010010000001000000110101010010110000111;
  c[5] = 132'b11000000100001100010000100000001001010000001010100100100110011011000011000011001100110001000010000000110111000000101001010010001100;
  c[6] = 132'b00110100000011110000000011000000101111101000000001100101000100100011100110111000000100101001100000000000100100000000100100001000000;
  c[7] = 132'b01110000100000001100000000000010101111000000001011000010101100100000111110110000010101100110100011000000000110100000100100010000110;
end

always@(posedge clock)
  if(clock == 1'b1 & k <8)
  begin
    Aout = c[k][63:0];
    Bout = c[k][127:64];
    op = c[k][131:128];
    k = k + 1;
  end
  else if(clock == 1'b0)
  begin
    d[k] = Din;
  end

endmodule
